
module System (
	clk_clk);	

	input		clk_clk;
endmodule
