
module System (
	clk_clk,
	uart_0_external_connection_rxd,
	uart_0_external_connection_txd);	

	input		clk_clk;
	input		uart_0_external_connection_rxd;
	output		uart_0_external_connection_txd;
endmodule
