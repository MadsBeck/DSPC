package BlockDecomp is
        type StringText is array(63 downto 0) of bit_vector(31 downto 0);
		type Constant_k is array(63 downto 0) of bit_vector(31 downto 0);
		type InitH is array (7 downto 0) of bit_vector(31 downto 0);
		
		
		constant Hcon : InitH := (
		X"6a09e667", X"bb67ae85", X"3c6ef372",X"a54ff53a",
		X"510e527f", X"9b05688c",X"1f83d9ab", X"5be0cd19");
								   
		constant constants : Constant_k := (
			x"428a2f98", x"71374491", x"b5c0fbcf", x"e9b5dba5", x"3956c25b", x"59f111f1", x"923f82a4", x"ab1c5ed5",
			x"d807aa98", x"12835b01", x"243185be", x"550c7dc3", x"72be5d74", x"80deb1fe", x"9bdc06a7", x"c19bf174",
			x"e49b69c1", x"efbe4786", x"0fc19dc6", x"240ca1cc", x"2de92c6f", x"4a7484aa", x"5cb0a9dc", x"76f988da",
			x"983e5152", x"a831c66d", x"b00327c8", x"bf597fc7", x"c6e00bf3", x"d5a79147", x"06ca6351", x"14292967",
			x"27b70a85", x"2e1b2138", x"4d2c6dfc", x"53380d13", x"650a7354", x"766a0abb", x"81c2c92e", x"92722c85",
			x"a2bfe8a1", x"a81a664b", x"c24b8b70", x"c76c51a3", x"d192e819", x"d6990624", x"f40e3585", x"106aa070",
			x"19a4c116", x"1e376c08", x"2748774c", x"34b0bcb5", x"391c0cb3", x"4ed8aa4a", x"5b9cca4f", x"682e6ff3",
			x"748f82ee", x"78a5636f", x"84c87814", x"8cc70208", x"90befffa", x"a4506ceb", x"bef9a3f7", x"c67178f2"
		);
		
end package;






entity HashComp is
	port(
		clk    : in std_logic;
		reset  : in std_logic;

		ready  : out std_logic; -- Ready to process the next block
		newData : in  std_logic; -- Start processing the next 
		
		input : IN StringText;
		output : OUT bit_vector(255 downto 0);

	);
end entity HashComp;


architecture rtl of HashComp is

	state_type is (IDLE,BUSY,DONE)
	signal state : state_type;
	
	signal h0, h1, h2, h3, h4, h5, h6, h7 : bit_vector(31 downto 0);
	
	signal T1, T2, a, b, c, d, e, f, g, h : bit_vector(31 downto 0);
	



begin

	output <= h0 & h1 & h2 & h3 & h4 & h5 & h6 & h7;
	
	ready <= '1' when state = IDLE else '0';
	
	
	   ---------------------------------------------------------------------------------------------------
   --! HashComp process
   ---------------------------------------------------------------------------------------------------
   hashCompProc : process(rst, clk)
   begin
      if (reset = '1') then
		a <= InitH(0);
		b <= InitH(1);
		c <= InitH(2);
		d <= InitH(3);
		e <= InitH(4);
		f <= InitH(5);
		g <= InitH(6);
		h <= InitH(7);
		T1 <= (others => '0');
		T2 <= (others => '0');
		
		state <= IDLE;
		

      elsif (clk'event and clk = '1') then
	  case state is
		when IDLE =>
			if (newData = '1') then
				
				state <= BUSY;
				
			end if;
		when BUSY =>
			for I 0 to 63 loop
			
			
			
			end loop;
				
	  
	  
	  

      end if;
   end process;

	








end architecture rtl;